** Profile: "SCHEMATIC1-bias"  [ c:\users\ddurachk\desktop\projects\grams\2 - schematics and layouts\100 - gse\simulation_folder\stability\lc_circuit-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\ddurachk\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "$(GRAMS)\PARTS\ISL70417SEH\isl70417.lib" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 20 10 10G
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
